
module REG100( clk, data, reset, enSig, outSig, outData );
  input [15:0] data;
  input [5:0] enSig;
  input [5:0] outSig;
  output [15:0] outData;
  input clk, reset;
  wire   N101, N102, N104, N105, N107, N108, N111, N113, N114, N116, N117,
         N120, N122, N123, N125, N126, N128, N129, N131, N132, N134, N135,
         N137, N138, N140, N141, N143, N144, N147, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n182, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n210, n211, n212, n213, n214, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n234, n235, n237, n238, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470;
  wire   [15:0] reg3;
  wire   [15:0] reg2;
  wire   [15:0] reg1;
  wire   [15:0] reg0;
  tri   [15:0] outData;

  DFFX2 \outData_tri_enable_reg[15]  ( .D(n411), .CLK(clk), .Q(N102), .QN(n204) );
  DFFX2 \outData_tri_enable_reg[14]  ( .D(n410), .CLK(clk), .Q(N105), .QN(n206) );
  DFFX2 \outData_tri_enable_reg[13]  ( .D(n409), .CLK(clk), .Q(N108), .QN(n208) );
  DFFX2 \outData_tri_enable_reg[12]  ( .D(n408), .CLK(clk), .Q(N111), .QN(n210) );
  DFFX2 \outData_tri_enable_reg[11]  ( .D(n407), .CLK(clk), .Q(N114), .QN(n212) );
  DFFX2 \outData_tri_enable_reg[10]  ( .D(n406), .CLK(clk), .Q(N117), .QN(n214) );
  DFFX2 \outData_tri_enable_reg[9]  ( .D(n405), .CLK(clk), .Q(N120), .QN(n216)
         );
  DFFX2 \outData_tri_enable_reg[8]  ( .D(n404), .CLK(clk), .Q(N123), .QN(n218)
         );
  DFFX2 \outData_tri_enable_reg[7]  ( .D(n403), .CLK(clk), .Q(N126), .QN(n220)
         );
  DFFX2 \outData_tri_enable_reg[6]  ( .D(n402), .CLK(clk), .Q(N129), .QN(n222)
         );
  DFFX2 \outData_tri_enable_reg[5]  ( .D(n401), .CLK(clk), .Q(N132), .QN(n224)
         );
  DFFX2 \outData_tri_enable_reg[4]  ( .D(n400), .CLK(clk), .Q(N135), .QN(n226)
         );
  DFFX2 \outData_tri_enable_reg[3]  ( .D(n399), .CLK(clk), .Q(N138), .QN(n228)
         );
  DFFX2 \outData_tri_enable_reg[2]  ( .D(n398), .CLK(clk), .Q(N141), .QN(n230)
         );
  DFFX2 \outData_tri_enable_reg[1]  ( .D(n397), .CLK(clk), .Q(N144), .QN(n232)
         );
  DFFX2 \outData_tri_enable_reg[0]  ( .D(n396), .CLK(clk), .Q(N147), .QN(n234)
         );
  DFFARX2 \reg2_reg[15]  ( .D(n395), .CLK(clk), .RSTB(n462), .Q(reg2[15]), 
        .QN(n290) );
  DFFARX2 \reg2_reg[14]  ( .D(n394), .CLK(clk), .RSTB(n466), .Q(reg2[14]), 
        .QN(n289) );
  DFFARX2 \reg2_reg[13]  ( .D(n393), .CLK(clk), .RSTB(n470), .Q(reg2[13]), 
        .QN(n288) );
  DFFARX2 \reg2_reg[12]  ( .D(n392), .CLK(clk), .RSTB(n466), .Q(reg2[12]), 
        .QN(n287) );
  DFFARX2 \reg2_reg[11]  ( .D(n391), .CLK(clk), .RSTB(n463), .Q(reg2[11]), 
        .QN(n286) );
  DFFARX2 \reg2_reg[10]  ( .D(n390), .CLK(clk), .RSTB(n466), .Q(reg2[10]), 
        .QN(n285) );
  DFFARX2 \reg2_reg[9]  ( .D(n389), .CLK(clk), .RSTB(n465), .Q(reg2[9]), .QN(
        n299) );
  DFFARX2 \reg2_reg[8]  ( .D(n388), .CLK(clk), .RSTB(n461), .Q(reg2[8]), .QN(
        n298) );
  DFFARX2 \reg2_reg[7]  ( .D(n387), .CLK(clk), .RSTB(n466), .Q(reg2[7]), .QN(
        n297) );
  DFFARX2 \reg2_reg[6]  ( .D(n386), .CLK(clk), .RSTB(n470), .Q(reg2[6]), .QN(
        n296) );
  DFFARX2 \reg2_reg[5]  ( .D(n385), .CLK(clk), .RSTB(n466), .Q(reg2[5]), .QN(
        n295) );
  DFFARX2 \reg2_reg[4]  ( .D(n384), .CLK(clk), .RSTB(n469), .Q(reg2[4]), .QN(
        n294) );
  DFFARX2 \reg2_reg[3]  ( .D(n383), .CLK(clk), .RSTB(n466), .Q(reg2[3]), .QN(
        n293) );
  DFFARX2 \reg2_reg[2]  ( .D(n382), .CLK(clk), .RSTB(n462), .Q(reg2[2]), .QN(
        n292) );
  DFFARX2 \reg2_reg[1]  ( .D(n381), .CLK(clk), .RSTB(n466), .Q(reg2[1]), .QN(
        n291) );
  DFFARX2 \reg2_reg[0]  ( .D(n380), .CLK(clk), .RSTB(n463), .Q(reg2[0]), .QN(
        n284) );
  DFFARX2 \reg1_reg[15]  ( .D(n379), .CLK(clk), .RSTB(n470), .Q(reg1[15]), 
        .QN(n274) );
  DFFARX2 \reg1_reg[14]  ( .D(n378), .CLK(clk), .RSTB(n467), .Q(reg1[14]), 
        .QN(n273) );
  DFFARX2 \reg1_reg[13]  ( .D(n377), .CLK(clk), .RSTB(n469), .Q(reg1[13]), 
        .QN(n272) );
  DFFARX2 \reg1_reg[12]  ( .D(n376), .CLK(clk), .RSTB(n467), .Q(reg1[12]), 
        .QN(n271) );
  DFFARX2 \reg1_reg[11]  ( .D(n375), .CLK(clk), .RSTB(n468), .Q(reg1[11]), 
        .QN(n270) );
  DFFARX2 \reg1_reg[10]  ( .D(n374), .CLK(clk), .RSTB(n467), .Q(reg1[10]), 
        .QN(n269) );
  DFFARX2 \reg1_reg[9]  ( .D(n373), .CLK(clk), .RSTB(n466), .Q(reg1[9]), .QN(
        n283) );
  DFFARX2 \reg1_reg[8]  ( .D(n372), .CLK(clk), .RSTB(n470), .Q(reg1[8]), .QN(
        n282) );
  DFFARX2 \reg1_reg[7]  ( .D(n371), .CLK(clk), .RSTB(n466), .Q(reg1[7]), .QN(
        n281) );
  DFFARX2 \reg1_reg[6]  ( .D(n370), .CLK(clk), .RSTB(n469), .Q(reg1[6]), .QN(
        n280) );
  DFFARX2 \reg1_reg[5]  ( .D(n369), .CLK(clk), .RSTB(n467), .Q(reg1[5]), .QN(
        n279) );
  DFFARX2 \reg1_reg[4]  ( .D(n368), .CLK(clk), .RSTB(n470), .Q(reg1[4]), .QN(
        n278) );
  DFFARX2 \reg1_reg[3]  ( .D(n367), .CLK(clk), .RSTB(n467), .Q(reg1[3]), .QN(
        n277) );
  DFFARX2 \reg1_reg[2]  ( .D(n366), .CLK(clk), .RSTB(n468), .Q(reg1[2]), .QN(
        n276) );
  DFFARX2 \reg1_reg[1]  ( .D(n365), .CLK(clk), .RSTB(n467), .Q(reg1[1]), .QN(
        n275) );
  DFFARX2 \reg1_reg[0]  ( .D(n364), .CLK(clk), .RSTB(n470), .Q(reg1[0]), .QN(
        n268) );
  DFFARX2 \reg0_reg[15]  ( .D(n363), .CLK(clk), .RSTB(n468), .Q(reg0[15]), 
        .QN(n258) );
  DFFARX2 \reg0_reg[14]  ( .D(n362), .CLK(clk), .RSTB(n468), .Q(reg0[14]), 
        .QN(n257) );
  DFFARX2 \reg0_reg[13]  ( .D(n361), .CLK(clk), .RSTB(n469), .Q(reg0[13]), 
        .QN(n256) );
  DFFARX2 \reg0_reg[12]  ( .D(n360), .CLK(clk), .RSTB(n468), .Q(reg0[12]), 
        .QN(n255) );
  DFFARX2 \reg0_reg[11]  ( .D(n359), .CLK(clk), .RSTB(n469), .Q(reg0[11]), 
        .QN(n254) );
  DFFARX2 \reg0_reg[10]  ( .D(n358), .CLK(clk), .RSTB(n468), .Q(reg0[10]), 
        .QN(n253) );
  DFFARX2 \reg0_reg[9]  ( .D(n357), .CLK(clk), .RSTB(n467), .Q(reg0[9]), .QN(
        n267) );
  DFFARX2 \reg0_reg[8]  ( .D(n356), .CLK(clk), .RSTB(n470), .Q(reg0[8]), .QN(
        n266) );
  DFFARX2 \reg0_reg[7]  ( .D(n355), .CLK(clk), .RSTB(n467), .Q(reg0[7]), .QN(
        n265) );
  DFFARX2 \reg0_reg[6]  ( .D(n354), .CLK(clk), .RSTB(n469), .Q(reg0[6]), .QN(
        n264) );
  DFFARX2 \reg0_reg[5]  ( .D(n353), .CLK(clk), .RSTB(n467), .Q(reg0[5]), .QN(
        n263) );
  DFFARX2 \reg0_reg[4]  ( .D(n352), .CLK(clk), .RSTB(n469), .Q(reg0[4]), .QN(
        n262) );
  DFFARX2 \reg0_reg[3]  ( .D(n351), .CLK(clk), .RSTB(n468), .Q(reg0[3]), .QN(
        n261) );
  DFFARX2 \reg0_reg[2]  ( .D(n350), .CLK(clk), .RSTB(n469), .Q(reg0[2]), .QN(
        n260) );
  DFFARX2 \reg0_reg[1]  ( .D(n349), .CLK(clk), .RSTB(n468), .Q(reg0[1]), .QN(
        n259) );
  DFFARX2 \reg0_reg[0]  ( .D(n348), .CLK(clk), .RSTB(n469), .Q(reg0[0]), .QN(
        n252) );
  DFFARX2 \reg3_reg[15]  ( .D(n347), .CLK(clk), .RSTB(n461), .Q(reg3[15]), 
        .QN(n306) );
  DFFX2 \outData_reg[15]  ( .D(n346), .CLK(clk), .Q(N101), .QN(n242) );
  DFFARX2 \reg3_reg[14]  ( .D(n345), .CLK(clk), .RSTB(n465), .Q(reg3[14]), 
        .QN(n305) );
  DFFX2 \outData_reg[14]  ( .D(n344), .CLK(clk), .Q(N104), .QN(n241) );
  DFFARX2 \reg3_reg[13]  ( .D(n343), .CLK(clk), .RSTB(n470), .Q(reg3[13]), 
        .QN(n304) );
  DFFX2 \outData_reg[13]  ( .D(n342), .CLK(clk), .Q(N107), .QN(n240) );
  DFFARX2 \reg3_reg[12]  ( .D(n341), .CLK(clk), .RSTB(n465), .Q(reg3[12]), 
        .QN(n303) );
  DFFX2 \outData_reg[12]  ( .D(n340), .CLK(clk), .Q(n416) );
  DFFARX2 \reg3_reg[11]  ( .D(n339), .CLK(clk), .RSTB(n462), .Q(reg3[11]), 
        .QN(n302) );
  DFFX2 \outData_reg[11]  ( .D(n338), .CLK(clk), .Q(N113), .QN(n238) );
  DFFARX2 \reg3_reg[10]  ( .D(n337), .CLK(clk), .RSTB(n465), .Q(reg3[10]), 
        .QN(n301) );
  DFFX2 \outData_reg[10]  ( .D(n336), .CLK(clk), .Q(N116), .QN(n237) );
  DFFARX2 \reg3_reg[9]  ( .D(n335), .CLK(clk), .RSTB(n468), .Q(reg3[9]), .QN(
        n315) );
  DFFX2 \outData_reg[9]  ( .D(n334), .CLK(clk), .Q(n417) );
  DFFARX2 \reg3_reg[8]  ( .D(n333), .CLK(clk), .RSTB(n465), .Q(reg3[8]), .QN(
        n314) );
  DFFX2 \outData_reg[8]  ( .D(n332), .CLK(clk), .Q(N122), .QN(n250) );
  DFFARX2 \reg3_reg[7]  ( .D(n331), .CLK(clk), .RSTB(n465), .Q(reg3[7]), .QN(
        n313) );
  DFFX2 \outData_reg[7]  ( .D(n330), .CLK(clk), .Q(N125), .QN(n249) );
  DFFARX2 \reg3_reg[6]  ( .D(n329), .CLK(clk), .RSTB(n470), .Q(reg3[6]), .QN(
        n312) );
  DFFX2 \outData_reg[6]  ( .D(n328), .CLK(clk), .Q(N128), .QN(n248) );
  DFFARX2 \reg3_reg[5]  ( .D(n327), .CLK(clk), .RSTB(n465), .Q(reg3[5]), .QN(
        n311) );
  DFFX2 \outData_reg[5]  ( .D(n326), .CLK(clk), .Q(N131), .QN(n247) );
  DFFARX2 \reg3_reg[4]  ( .D(n325), .CLK(clk), .RSTB(n462), .Q(reg3[4]), .QN(
        n310) );
  DFFX2 \outData_reg[4]  ( .D(n324), .CLK(clk), .Q(N134), .QN(n246) );
  DFFARX2 \reg3_reg[3]  ( .D(n323), .CLK(clk), .RSTB(n465), .Q(reg3[3]), .QN(
        n309) );
  DFFX2 \outData_reg[3]  ( .D(n322), .CLK(clk), .Q(N137), .QN(n245) );
  DFFARX2 \reg3_reg[2]  ( .D(n321), .CLK(clk), .RSTB(n463), .Q(reg3[2]), .QN(
        n308) );
  DFFX2 \outData_reg[2]  ( .D(n320), .CLK(clk), .Q(N140), .QN(n244) );
  DFFARX2 \reg3_reg[1]  ( .D(n319), .CLK(clk), .RSTB(n465), .Q(reg3[1]), .QN(
        n307) );
  DFFX2 \outData_reg[1]  ( .D(n318), .CLK(clk), .Q(N143), .QN(n243) );
  DFFARX2 \reg3_reg[0]  ( .D(n317), .CLK(clk), .RSTB(n461), .Q(reg3[0]), .QN(
        n300) );
  DFFX2 \outData_reg[0]  ( .D(n316), .CLK(clk), .Q(n418) );
  TNBUFFHX8 \outData_tri[0]  ( .IN(n441), .ENB(n434), .Q(outData[0]) );
  TNBUFFHX8 \outData_tri[1]  ( .IN(n438), .ENB(n433), .Q(outData[1]) );
  TNBUFFHX8 \outData_tri[2]  ( .IN(n442), .ENB(n432), .Q(outData[2]) );
  TNBUFFHX8 \outData_tri[3]  ( .IN(n435), .ENB(n431), .Q(outData[3]) );
  TNBUFFHX8 \outData_tri[4]  ( .IN(n447), .ENB(n430), .Q(outData[4]) );
  TNBUFFHX8 \outData_tri[5]  ( .IN(n439), .ENB(n429), .Q(outData[5]) );
  TNBUFFHX8 \outData_tri[6]  ( .IN(n449), .ENB(n428), .Q(outData[6]) );
  TNBUFFHX8 \outData_tri[7]  ( .IN(n440), .ENB(n427), .Q(outData[7]) );
  TNBUFFHX8 \outData_tri[8]  ( .IN(n443), .ENB(n426), .Q(outData[8]) );
  TNBUFFHX8 \outData_tri[9]  ( .IN(n436), .ENB(n425), .Q(outData[9]) );
  TNBUFFHX8 \outData_tri[10]  ( .IN(n437), .ENB(n424), .Q(outData[10]) );
  TNBUFFHX8 \outData_tri[11]  ( .IN(n444), .ENB(n423), .Q(outData[11]) );
  TNBUFFHX8 \outData_tri[12]  ( .IN(n445), .ENB(n422), .Q(outData[12]) );
  TNBUFFHX8 \outData_tri[13]  ( .IN(n448), .ENB(n421), .Q(outData[13]) );
  TNBUFFHX8 \outData_tri[14]  ( .IN(n450), .ENB(n420), .Q(outData[14]) );
  TNBUFFHX8 \outData_tri[15]  ( .IN(n446), .ENB(n419), .Q(outData[15]) );
  AO22X2 U2 ( .IN1(data[9]), .IN2(n460), .IN3(n459), .IN4(n83), .Q(n335) );
  AO22X2 U3 ( .IN1(data[8]), .IN2(n460), .IN3(n459), .IN4(n84), .Q(n333) );
  AO22X2 U4 ( .IN1(data[7]), .IN2(n460), .IN3(n459), .IN4(n85), .Q(n331) );
  AO22X2 U5 ( .IN1(data[6]), .IN2(n460), .IN3(n459), .IN4(n86), .Q(n329) );
  AO22X2 U6 ( .IN1(data[5]), .IN2(n460), .IN3(n459), .IN4(n87), .Q(n327) );
  AO22X2 U7 ( .IN1(data[4]), .IN2(n460), .IN3(n459), .IN4(n88), .Q(n325) );
  AO22X2 U8 ( .IN1(data[3]), .IN2(n460), .IN3(n459), .IN4(n89), .Q(n323) );
  AO22X2 U9 ( .IN1(data[2]), .IN2(n460), .IN3(n459), .IN4(n90), .Q(n321) );
  AO22X2 U10 ( .IN1(data[1]), .IN2(n460), .IN3(n459), .IN4(n91), .Q(n319) );
  AO22X2 U11 ( .IN1(data[15]), .IN2(n460), .IN3(n459), .IN4(n92), .Q(n347) );
  AO22X2 U12 ( .IN1(data[14]), .IN2(n460), .IN3(n459), .IN4(n93), .Q(n345) );
  AO22X2 U13 ( .IN1(data[13]), .IN2(n460), .IN3(n459), .IN4(n94), .Q(n343) );
  AO22X2 U14 ( .IN1(data[12]), .IN2(n460), .IN3(n459), .IN4(n95), .Q(n341) );
  AO22X2 U15 ( .IN1(data[11]), .IN2(n460), .IN3(n459), .IN4(n96), .Q(n339) );
  AO22X2 U16 ( .IN1(data[10]), .IN2(n460), .IN3(n459), .IN4(n97), .Q(n337) );
  AO22X2 U17 ( .IN1(data[0]), .IN2(n460), .IN3(n459), .IN4(n98), .Q(n317) );
  NAND4X0 U19 ( .IN1(enSig[2]), .IN2(enSig[1]), .IN3(enSig[0]), .IN4(n99), 
        .QN(n82) );
  AO22X2 U20 ( .IN1(n458), .IN2(data[9]), .IN3(n457), .IN4(n102), .Q(n389) );
  AO22X2 U21 ( .IN1(n458), .IN2(data[8]), .IN3(n457), .IN4(n103), .Q(n388) );
  AO22X2 U22 ( .IN1(n458), .IN2(data[7]), .IN3(n457), .IN4(n104), .Q(n387) );
  AO22X2 U23 ( .IN1(n458), .IN2(data[6]), .IN3(n457), .IN4(n105), .Q(n386) );
  AO22X2 U24 ( .IN1(n458), .IN2(data[5]), .IN3(n457), .IN4(n106), .Q(n385) );
  AO22X2 U25 ( .IN1(n458), .IN2(data[4]), .IN3(n457), .IN4(n107), .Q(n384) );
  AO22X2 U26 ( .IN1(n458), .IN2(data[3]), .IN3(n457), .IN4(n108), .Q(n383) );
  AO22X2 U27 ( .IN1(n458), .IN2(data[2]), .IN3(n457), .IN4(n109), .Q(n382) );
  AO22X2 U28 ( .IN1(n458), .IN2(data[1]), .IN3(n457), .IN4(n110), .Q(n381) );
  AO22X2 U29 ( .IN1(n458), .IN2(data[15]), .IN3(n457), .IN4(n111), .Q(n395) );
  AO22X2 U30 ( .IN1(n458), .IN2(data[14]), .IN3(n457), .IN4(n112), .Q(n394) );
  AO22X2 U31 ( .IN1(n458), .IN2(data[13]), .IN3(n457), .IN4(n113), .Q(n393) );
  AO22X2 U32 ( .IN1(n458), .IN2(data[12]), .IN3(n457), .IN4(n114), .Q(n392) );
  AO22X2 U33 ( .IN1(n458), .IN2(data[11]), .IN3(n457), .IN4(n115), .Q(n391) );
  AO22X2 U34 ( .IN1(n458), .IN2(data[10]), .IN3(n457), .IN4(n116), .Q(n390) );
  AO22X2 U35 ( .IN1(n458), .IN2(data[0]), .IN3(n457), .IN4(n117), .Q(n380) );
  NAND3X0 U37 ( .IN1(enSig[1]), .IN2(enSig[0]), .IN3(n118), .QN(n101) );
  AO22X2 U38 ( .IN1(n456), .IN2(data[9]), .IN3(n455), .IN4(n121), .Q(n373) );
  AO22X2 U39 ( .IN1(n456), .IN2(data[8]), .IN3(n455), .IN4(n122), .Q(n372) );
  AO22X2 U40 ( .IN1(n456), .IN2(data[7]), .IN3(n455), .IN4(n123), .Q(n371) );
  AO22X2 U41 ( .IN1(n456), .IN2(data[6]), .IN3(n455), .IN4(n124), .Q(n370) );
  AO22X2 U42 ( .IN1(n456), .IN2(data[5]), .IN3(n455), .IN4(n125), .Q(n369) );
  AO22X2 U43 ( .IN1(n456), .IN2(data[4]), .IN3(n455), .IN4(n126), .Q(n368) );
  AO22X2 U44 ( .IN1(n456), .IN2(data[3]), .IN3(n455), .IN4(n127), .Q(n367) );
  AO22X2 U45 ( .IN1(n456), .IN2(data[2]), .IN3(n455), .IN4(n128), .Q(n366) );
  AO22X2 U46 ( .IN1(n456), .IN2(data[1]), .IN3(n455), .IN4(n129), .Q(n365) );
  AO22X2 U47 ( .IN1(n456), .IN2(data[15]), .IN3(n455), .IN4(n130), .Q(n379) );
  AO22X2 U48 ( .IN1(n456), .IN2(data[14]), .IN3(n455), .IN4(n131), .Q(n378) );
  AO22X2 U49 ( .IN1(n456), .IN2(data[13]), .IN3(n455), .IN4(n132), .Q(n377) );
  AO22X2 U50 ( .IN1(n456), .IN2(data[12]), .IN3(n455), .IN4(n133), .Q(n376) );
  AO22X2 U51 ( .IN1(n456), .IN2(data[11]), .IN3(n455), .IN4(n134), .Q(n375) );
  AO22X2 U52 ( .IN1(n456), .IN2(data[10]), .IN3(n455), .IN4(n135), .Q(n374) );
  AO22X2 U53 ( .IN1(n456), .IN2(data[0]), .IN3(n455), .IN4(n136), .Q(n364) );
  NAND3X0 U55 ( .IN1(enSig[0]), .IN2(n137), .IN3(n118), .QN(n120) );
  AO22X2 U56 ( .IN1(n454), .IN2(data[9]), .IN3(n453), .IN4(n140), .Q(n357) );
  AO22X2 U57 ( .IN1(n454), .IN2(data[8]), .IN3(n453), .IN4(n141), .Q(n356) );
  AO22X2 U58 ( .IN1(n454), .IN2(data[7]), .IN3(n453), .IN4(n142), .Q(n355) );
  AO22X2 U59 ( .IN1(n454), .IN2(data[6]), .IN3(n453), .IN4(n143), .Q(n354) );
  AO22X2 U60 ( .IN1(n454), .IN2(data[5]), .IN3(n453), .IN4(n144), .Q(n353) );
  AO22X2 U61 ( .IN1(n454), .IN2(data[4]), .IN3(n453), .IN4(n145), .Q(n352) );
  AO22X2 U62 ( .IN1(n454), .IN2(data[3]), .IN3(n453), .IN4(n146), .Q(n351) );
  AO22X2 U63 ( .IN1(n454), .IN2(data[2]), .IN3(n453), .IN4(n147), .Q(n350) );
  AO22X2 U64 ( .IN1(n454), .IN2(data[1]), .IN3(n453), .IN4(n148), .Q(n349) );
  AO22X2 U65 ( .IN1(n454), .IN2(data[15]), .IN3(n453), .IN4(n149), .Q(n363) );
  AO22X2 U66 ( .IN1(n454), .IN2(data[14]), .IN3(n453), .IN4(n150), .Q(n362) );
  AO22X2 U67 ( .IN1(n454), .IN2(data[13]), .IN3(n453), .IN4(n151), .Q(n361) );
  AO22X2 U68 ( .IN1(n454), .IN2(data[12]), .IN3(n453), .IN4(n152), .Q(n360) );
  AO22X2 U69 ( .IN1(n454), .IN2(data[11]), .IN3(n453), .IN4(n153), .Q(n359) );
  AO22X2 U70 ( .IN1(n454), .IN2(data[10]), .IN3(n453), .IN4(n154), .Q(n358) );
  AO22X2 U71 ( .IN1(n454), .IN2(data[0]), .IN3(n453), .IN4(n155), .Q(n348) );
  NAND3X0 U73 ( .IN1(n156), .IN2(n137), .IN3(n118), .QN(n139) );
  ISOLANDX1 U74 ( .D(n99), .ISO(enSig[2]), .Q(n118) );
  NOR3X0 U75 ( .IN1(enSig[5]), .IN2(enSig[4]), .IN3(enSig[3]), .QN(n99) );
  NAND2X0 U78 ( .IN1(n157), .IN2(n158), .QN(n405) );
  NAND2X0 U80 ( .IN1(n157), .IN2(n159), .QN(n404) );
  NAND2X0 U82 ( .IN1(n157), .IN2(n160), .QN(n403) );
  NAND2X0 U84 ( .IN1(n157), .IN2(n161), .QN(n402) );
  NAND2X0 U86 ( .IN1(n157), .IN2(n162), .QN(n401) );
  NAND2X0 U88 ( .IN1(n157), .IN2(n163), .QN(n400) );
  NAND2X0 U90 ( .IN1(n157), .IN2(n164), .QN(n399) );
  NAND2X0 U92 ( .IN1(n157), .IN2(n165), .QN(n398) );
  NAND2X0 U94 ( .IN1(n157), .IN2(n166), .QN(n397) );
  NAND2X0 U96 ( .IN1(n157), .IN2(n167), .QN(n411) );
  NAND2X0 U98 ( .IN1(n157), .IN2(n168), .QN(n410) );
  NAND2X0 U100 ( .IN1(n157), .IN2(n169), .QN(n409) );
  NAND2X0 U102 ( .IN1(n157), .IN2(n170), .QN(n408) );
  NAND2X0 U104 ( .IN1(n157), .IN2(n171), .QN(n407) );
  NAND2X0 U106 ( .IN1(n157), .IN2(n172), .QN(n406) );
  NAND2X0 U108 ( .IN1(n157), .IN2(n173), .QN(n396) );
  NOR2X1 U112 ( .IN1(reset), .IN2(n178), .QN(n176) );
  AO221X2 U113 ( .IN1(n179), .IN2(n102), .IN3(reset), .IN4(n436), .IN5(n180), 
        .Q(n334) );
  AO222X2 U114 ( .IN1(n451), .IN2(n140), .IN3(n182), .IN4(n83), .IN5(n452), 
        .IN6(n121), .Q(n180) );
  AO221X2 U120 ( .IN1(n179), .IN2(n103), .IN3(reset), .IN4(n443), .IN5(n184), 
        .Q(n332) );
  AO222X2 U121 ( .IN1(n451), .IN2(n141), .IN3(n182), .IN4(n84), .IN5(n452), 
        .IN6(n122), .Q(n184) );
  AO221X2 U127 ( .IN1(n179), .IN2(n104), .IN3(reset), .IN4(n440), .IN5(n185), 
        .Q(n330) );
  AO222X2 U128 ( .IN1(n451), .IN2(n142), .IN3(n182), .IN4(n85), .IN5(n452), 
        .IN6(n123), .Q(n185) );
  AO221X2 U134 ( .IN1(n179), .IN2(n105), .IN3(reset), .IN4(n449), .IN5(n186), 
        .Q(n328) );
  AO222X2 U135 ( .IN1(n451), .IN2(n143), .IN3(n182), .IN4(n86), .IN5(n452), 
        .IN6(n124), .Q(n186) );
  AO221X2 U141 ( .IN1(n179), .IN2(n106), .IN3(reset), .IN4(n439), .IN5(n187), 
        .Q(n326) );
  AO222X2 U142 ( .IN1(n451), .IN2(n144), .IN3(n182), .IN4(n87), .IN5(n452), 
        .IN6(n125), .Q(n187) );
  AO221X2 U148 ( .IN1(n179), .IN2(n107), .IN3(reset), .IN4(n447), .IN5(n188), 
        .Q(n324) );
  AO222X2 U149 ( .IN1(n451), .IN2(n145), .IN3(n182), .IN4(n88), .IN5(n452), 
        .IN6(n126), .Q(n188) );
  AO221X2 U155 ( .IN1(n179), .IN2(n108), .IN3(reset), .IN4(n435), .IN5(n189), 
        .Q(n322) );
  AO222X2 U156 ( .IN1(n451), .IN2(n146), .IN3(n182), .IN4(n89), .IN5(n452), 
        .IN6(n127), .Q(n189) );
  AO221X2 U162 ( .IN1(n179), .IN2(n109), .IN3(reset), .IN4(n442), .IN5(n190), 
        .Q(n320) );
  AO222X2 U163 ( .IN1(n451), .IN2(n147), .IN3(n182), .IN4(n90), .IN5(n452), 
        .IN6(n128), .Q(n190) );
  AO221X2 U169 ( .IN1(n179), .IN2(n110), .IN3(reset), .IN4(n438), .IN5(n191), 
        .Q(n318) );
  AO222X2 U170 ( .IN1(n451), .IN2(n148), .IN3(n182), .IN4(n91), .IN5(n452), 
        .IN6(n129), .Q(n191) );
  AO221X2 U176 ( .IN1(n179), .IN2(n111), .IN3(reset), .IN4(n446), .IN5(n192), 
        .Q(n346) );
  AO222X2 U177 ( .IN1(n451), .IN2(n149), .IN3(n182), .IN4(n92), .IN5(n452), 
        .IN6(n130), .Q(n192) );
  AO221X2 U183 ( .IN1(n179), .IN2(n112), .IN3(reset), .IN4(n450), .IN5(n193), 
        .Q(n344) );
  AO222X2 U184 ( .IN1(n451), .IN2(n150), .IN3(n182), .IN4(n93), .IN5(n452), 
        .IN6(n131), .Q(n193) );
  AO221X2 U190 ( .IN1(n179), .IN2(n113), .IN3(reset), .IN4(n448), .IN5(n194), 
        .Q(n342) );
  AO222X2 U191 ( .IN1(n451), .IN2(n151), .IN3(n182), .IN4(n94), .IN5(n452), 
        .IN6(n132), .Q(n194) );
  AO221X2 U197 ( .IN1(n179), .IN2(n114), .IN3(reset), .IN4(n445), .IN5(n195), 
        .Q(n340) );
  AO222X2 U198 ( .IN1(n451), .IN2(n152), .IN3(n182), .IN4(n95), .IN5(n452), 
        .IN6(n133), .Q(n195) );
  AO221X2 U204 ( .IN1(n179), .IN2(n115), .IN3(reset), .IN4(n444), .IN5(n196), 
        .Q(n338) );
  AO222X2 U205 ( .IN1(n451), .IN2(n153), .IN3(n182), .IN4(n96), .IN5(n452), 
        .IN6(n134), .Q(n196) );
  AO221X2 U211 ( .IN1(n179), .IN2(n116), .IN3(reset), .IN4(n437), .IN5(n197), 
        .Q(n336) );
  AO222X2 U212 ( .IN1(n451), .IN2(n154), .IN3(n182), .IN4(n97), .IN5(n452), 
        .IN6(n135), .Q(n197) );
  AO221X2 U218 ( .IN1(n179), .IN2(n117), .IN3(reset), .IN4(n441), .IN5(n198), 
        .Q(n316) );
  AO222X2 U219 ( .IN1(n451), .IN2(n155), .IN3(n182), .IN4(n98), .IN5(n452), 
        .IN6(n136), .Q(n198) );
  NAND3X0 U222 ( .IN1(n199), .IN2(n200), .IN3(outSig[0]), .QN(n177) );
  NAND4X0 U225 ( .IN1(outSig[2]), .IN2(outSig[1]), .IN3(outSig[0]), .IN4(n201), 
        .QN(n174) );
  NAND3X0 U228 ( .IN1(n202), .IN2(n200), .IN3(n199), .QN(n175) );
  ISOLANDX1 U233 ( .D(n178), .ISO(reset), .Q(n179) );
  AND3X1 U234 ( .IN1(outSig[0]), .IN2(n199), .IN3(outSig[1]), .Q(n178) );
  ISOLANDX1 U235 ( .D(n201), .ISO(outSig[2]), .Q(n199) );
  NOR3X0 U236 ( .IN1(outSig[5]), .IN2(outSig[4]), .IN3(outSig[3]), .QN(n201)
         );
  ISOLORX2 U237 ( .D(n175), .ISO(reset), .Q(n412) );
  ISOLORX2 U238 ( .D(n177), .ISO(reset), .Q(n413) );
  ISOLORX2 U239 ( .D(n174), .ISO(reset), .Q(n414) );
  INVX0 U240 ( .IN(n414), .QN(n182) );
  AND4X1 U241 ( .IN1(n174), .IN2(n175), .IN3(n176), .IN4(n177), .Q(n415) );
  INVX0 U242 ( .IN(n415), .QN(n157) );
  ISOLORX2 U243 ( .D(n464), .ISO(n434), .Q(n173) );
  ISOLORX2 U244 ( .D(n464), .ISO(n433), .Q(n166) );
  ISOLORX2 U245 ( .D(n464), .ISO(n429), .Q(n162) );
  ISOLORX2 U246 ( .D(n464), .ISO(n425), .Q(n158) );
  ISOLORX2 U247 ( .D(n464), .ISO(n423), .Q(n171) );
  ISOLORX2 U248 ( .D(n464), .ISO(n422), .Q(n170) );
  ISOLORX2 U249 ( .D(n464), .ISO(n420), .Q(n168) );
  NBUFFX16 U250 ( .IN(n204), .Q(n419) );
  OR2X2 U251 ( .IN1(n235), .IN2(n419), .Q(n167) );
  NBUFFX16 U252 ( .IN(n206), .Q(n420) );
  NBUFFX16 U253 ( .IN(n208), .Q(n421) );
  OR2X2 U254 ( .IN1(n235), .IN2(n421), .Q(n169) );
  NBUFFX16 U255 ( .IN(n210), .Q(n422) );
  NBUFFX16 U256 ( .IN(n212), .Q(n423) );
  NBUFFX16 U257 ( .IN(n214), .Q(n424) );
  OR2X2 U258 ( .IN1(n235), .IN2(n424), .Q(n172) );
  NBUFFX16 U259 ( .IN(n216), .Q(n425) );
  NBUFFX16 U260 ( .IN(n218), .Q(n426) );
  OR2X2 U261 ( .IN1(n235), .IN2(n426), .Q(n159) );
  NBUFFX16 U262 ( .IN(n220), .Q(n427) );
  OR2X2 U263 ( .IN1(n235), .IN2(n427), .Q(n160) );
  NBUFFX16 U264 ( .IN(n222), .Q(n428) );
  OR2X2 U265 ( .IN1(n235), .IN2(n428), .Q(n161) );
  NBUFFX16 U266 ( .IN(n224), .Q(n429) );
  NBUFFX16 U267 ( .IN(n226), .Q(n430) );
  OR2X2 U268 ( .IN1(n235), .IN2(n430), .Q(n163) );
  NBUFFX16 U269 ( .IN(n228), .Q(n431) );
  OR2X2 U270 ( .IN1(n235), .IN2(n431), .Q(n164) );
  NBUFFX16 U271 ( .IN(n230), .Q(n432) );
  OR2X2 U272 ( .IN1(n235), .IN2(n432), .Q(n165) );
  NBUFFX16 U273 ( .IN(n232), .Q(n433) );
  NBUFFX16 U274 ( .IN(n234), .Q(n434) );
  NBUFFX16 U275 ( .IN(n227), .Q(n435) );
  AOINVX1 U276 ( .IN(n245), .QN(n227) );
  NBUFFX16 U277 ( .IN(n417), .Q(n436) );
  NBUFFX16 U278 ( .IN(n213), .Q(n437) );
  AOINVX1 U279 ( .IN(n237), .QN(n213) );
  NBUFFX16 U280 ( .IN(n231), .Q(n438) );
  AOINVX1 U281 ( .IN(n243), .QN(n231) );
  NBUFFX16 U282 ( .IN(n223), .Q(n439) );
  AOINVX1 U283 ( .IN(n247), .QN(n223) );
  NBUFFX16 U284 ( .IN(n219), .Q(n440) );
  AOINVX1 U285 ( .IN(n249), .QN(n219) );
  NBUFFX16 U286 ( .IN(n418), .Q(n441) );
  NBUFFX16 U287 ( .IN(n229), .Q(n442) );
  AOINVX1 U288 ( .IN(n244), .QN(n229) );
  NBUFFX16 U289 ( .IN(n217), .Q(n443) );
  AOINVX1 U290 ( .IN(n250), .QN(n217) );
  NBUFFX16 U291 ( .IN(n211), .Q(n444) );
  AOINVX1 U292 ( .IN(n238), .QN(n211) );
  NBUFFX16 U293 ( .IN(n416), .Q(n445) );
  NBUFFX16 U294 ( .IN(n203), .Q(n446) );
  AOINVX1 U295 ( .IN(n242), .QN(n203) );
  NBUFFX16 U296 ( .IN(n225), .Q(n447) );
  AOINVX1 U297 ( .IN(n246), .QN(n225) );
  NBUFFX16 U298 ( .IN(n207), .Q(n448) );
  AOINVX1 U299 ( .IN(n240), .QN(n207) );
  NBUFFX16 U300 ( .IN(n221), .Q(n449) );
  AOINVX1 U301 ( .IN(n248), .QN(n221) );
  NBUFFX16 U302 ( .IN(n205), .Q(n450) );
  AOINVX1 U303 ( .IN(n241), .QN(n205) );
  AOBUFX1 U304 ( .IN(n462), .Q(n468) );
  AOBUFX1 U305 ( .IN(n462), .Q(n467) );
  AOBUFX1 U306 ( .IN(n463), .Q(n469) );
  AOBUFX1 U307 ( .IN(n463), .Q(n470) );
  AOBUFX1 U308 ( .IN(n461), .Q(n465) );
  AOBUFX1 U309 ( .IN(n461), .Q(n466) );
  AOBUFX1 U310 ( .IN(n461), .Q(n462) );
  AOBUFX1 U311 ( .IN(n461), .Q(n463) );
  AOINVX2 U312 ( .IN(n82), .QN(n460) );
  AOINVX2 U313 ( .IN(n139), .QN(n454) );
  AOINVX2 U314 ( .IN(n120), .QN(n456) );
  AOINVX2 U315 ( .IN(n101), .QN(n458) );
  AOBUFX1 U316 ( .IN(n464), .Q(n461) );
  AOBUFX1 U317 ( .IN(n235), .Q(n464) );
  AOINVX1 U318 ( .IN(outSig[0]), .QN(n202) );
  AOINVX2 U319 ( .IN(n412), .QN(n451) );
  AOINVX1 U320 ( .IN(reset), .QN(n235) );
  AOBUFX1 U321 ( .IN(n82), .Q(n459) );
  AOINVX1 U322 ( .IN(outSig[1]), .QN(n200) );
  AOINVX1 U323 ( .IN(enSig[1]), .QN(n137) );
  AOINVX2 U324 ( .IN(n413), .QN(n452) );
  AOBUFX1 U325 ( .IN(n139), .Q(n453) );
  AOINVX1 U326 ( .IN(enSig[0]), .QN(n156) );
  AOBUFX1 U327 ( .IN(n120), .Q(n455) );
  AOBUFX1 U328 ( .IN(n101), .Q(n457) );
  AOINVX1 U329 ( .IN(n284), .QN(n117) );
  AOINVX1 U330 ( .IN(n291), .QN(n110) );
  AOINVX1 U331 ( .IN(n292), .QN(n109) );
  AOINVX1 U332 ( .IN(n293), .QN(n108) );
  AOINVX1 U333 ( .IN(n294), .QN(n107) );
  AOINVX1 U334 ( .IN(n295), .QN(n106) );
  AOINVX1 U335 ( .IN(n296), .QN(n105) );
  AOINVX1 U336 ( .IN(n297), .QN(n104) );
  AOINVX1 U337 ( .IN(n298), .QN(n103) );
  AOINVX1 U338 ( .IN(n299), .QN(n102) );
  AOINVX1 U339 ( .IN(n285), .QN(n116) );
  AOINVX1 U340 ( .IN(n286), .QN(n115) );
  AOINVX1 U341 ( .IN(n287), .QN(n114) );
  AOINVX1 U342 ( .IN(n288), .QN(n113) );
  AOINVX1 U343 ( .IN(n289), .QN(n112) );
  AOINVX1 U344 ( .IN(n290), .QN(n111) );
  AOINVX1 U345 ( .IN(n300), .QN(n98) );
  AOINVX1 U346 ( .IN(n307), .QN(n91) );
  AOINVX1 U347 ( .IN(n308), .QN(n90) );
  AOINVX1 U348 ( .IN(n309), .QN(n89) );
  AOINVX1 U349 ( .IN(n310), .QN(n88) );
  AOINVX1 U350 ( .IN(n311), .QN(n87) );
  AOINVX1 U351 ( .IN(n312), .QN(n86) );
  AOINVX1 U352 ( .IN(n313), .QN(n85) );
  AOINVX1 U353 ( .IN(n314), .QN(n84) );
  AOINVX1 U354 ( .IN(n315), .QN(n83) );
  AOINVX1 U355 ( .IN(n301), .QN(n97) );
  AOINVX1 U356 ( .IN(n302), .QN(n96) );
  AOINVX1 U357 ( .IN(n303), .QN(n95) );
  AOINVX1 U358 ( .IN(n304), .QN(n94) );
  AOINVX1 U359 ( .IN(n305), .QN(n93) );
  AOINVX1 U360 ( .IN(n306), .QN(n92) );
  AOINVX1 U361 ( .IN(n268), .QN(n136) );
  AOINVX1 U362 ( .IN(n275), .QN(n129) );
  AOINVX1 U363 ( .IN(n276), .QN(n128) );
  AOINVX1 U364 ( .IN(n277), .QN(n127) );
  AOINVX1 U365 ( .IN(n278), .QN(n126) );
  AOINVX1 U366 ( .IN(n279), .QN(n125) );
  AOINVX1 U367 ( .IN(n280), .QN(n124) );
  AOINVX1 U368 ( .IN(n281), .QN(n123) );
  AOINVX1 U369 ( .IN(n282), .QN(n122) );
  AOINVX1 U370 ( .IN(n283), .QN(n121) );
  AOINVX1 U371 ( .IN(n269), .QN(n135) );
  AOINVX1 U372 ( .IN(n270), .QN(n134) );
  AOINVX1 U373 ( .IN(n271), .QN(n133) );
  AOINVX1 U374 ( .IN(n272), .QN(n132) );
  AOINVX1 U375 ( .IN(n273), .QN(n131) );
  AOINVX1 U376 ( .IN(n274), .QN(n130) );
  AOINVX1 U377 ( .IN(n252), .QN(n155) );
  AOINVX1 U378 ( .IN(n259), .QN(n148) );
  AOINVX1 U379 ( .IN(n260), .QN(n147) );
  AOINVX1 U380 ( .IN(n261), .QN(n146) );
  AOINVX1 U381 ( .IN(n262), .QN(n145) );
  AOINVX1 U382 ( .IN(n263), .QN(n144) );
  AOINVX1 U383 ( .IN(n264), .QN(n143) );
  AOINVX1 U384 ( .IN(n265), .QN(n142) );
  AOINVX1 U385 ( .IN(n266), .QN(n141) );
  AOINVX1 U386 ( .IN(n267), .QN(n140) );
  AOINVX1 U387 ( .IN(n253), .QN(n154) );
  AOINVX1 U388 ( .IN(n254), .QN(n153) );
  AOINVX1 U389 ( .IN(n255), .QN(n152) );
  AOINVX1 U390 ( .IN(n256), .QN(n151) );
  AOINVX1 U391 ( .IN(n257), .QN(n150) );
  AOINVX1 U392 ( .IN(n258), .QN(n149) );
endmodule

